package apb_pkg;
  import uvm_pkg::*;

  typedef uvm_config_db#(virtual apb_if) uvm_config_db#(virtual apb_if);
  `include "uvm_macros.svh"

  `include "apb_packet.sv"
  `include "apb_monitor.sv"
  `include "apb_sequencer.sv"
  `include "apb_seqs.sv"
  `include "apb_driver.sv"
  `include "apb_agent.sv"
  `include "apb_env.sv"
endpackage : apb_pkg